module InstMem (
        input wire ce,                // 存储器使能信号
        input wire [31:0] addr,       // 取指地址
        output wire [31:0] data       // 输出指令数据
    );

    reg [31:0] mem [0:1023];      // 1024 个 32 位的存储单元

    initial begin
        mem[0] = 32'h340800FF; // ORI $8, $0, 0xFF
        mem[1] = 32'h3409FF00; // ORI $9, $0, 0xFF00

        mem[2] = 32'h300A00FF; // ANDI $10, $0, 0xFF
        mem[3] = 32'h300BFF00; // ANDI $11, $0, 0xFF00

        mem[4] = 32'h200C0001; // ADDI $12, $0, 1
        mem[5] = 32'h200DFFFF; // ADDI $13, $0, -1

        mem[6] = 32'h240E0002; // SUBI $14, $0, 2 (using pseudo-instruction: ADDI $14, $0, -2)
        mem[7] = 32'h240FFFFE; // SUBI $15, $0, -2

        mem[8] = 32'h3C100003; // LUI $16, 0x0003
        mem[9] = 32'h3C1100FF; // LUI $17, 0x00FF

        mem[10] = 32'h02124024; // AND $8, $16, $18
        mem[11] = 32'h02314824; // AND $9, $17, $19

        mem[12] = 32'h02125026; // XOR $10, $16, $18
        mem[13] = 32'h02315826; // XOR $11, $17, $19

        mem[14] = 32'h02126020; // ADD $12, $16, $18
        mem[15] = 32'h02316820; // ADD $13, $17, $19

        mem[16] = 32'h02127022; // SUB $14, $16, $18
        mem[17] = 32'h02317822; // SUB $15, $17, $19

        mem[18] = 32'h00104080; // SLL $8, $8, 2
        mem[19] = 32'h00104880; // SLL $9, $9, 2

        mem[20] = 32'h00105082; // SRL $10, $10, 2
        mem[21] = 32'h00105882; // SRL $11, $11, 2

        mem[22] = 32'h00106083; // SRA $12, $12, 2
        mem[23] = 32'h00106883; // SRA $13, $13, 2

        // 测试 BEQ (当 $16 和 $17 相等时跳转)
        mem[24] = 32'h12110001; // BEQ $16, $17, offset=1 (跳转到 mem[25])

        // 测试 BNE (当 $16 和 $17 不相等时跳转)
        mem[25] = 32'h16110001; // BNE $16, $17, offset=1 (跳转到 mem[26])

        // 设置寄存器值使得 BEQ 和 BNE 测试通过
        // BEQ 跳转
        mem[26] = 32'h34010000; // ORI $1, $0, 0x0000 (设置 $16 = $17)，BEQ 跳转成立
        mem[27] = 32'h3402FFFF; // ORI $2, $0, 0xFFFF

        // 测试 JAL (跳转到指定地址并保存返回地址)
        mem[28] = 32'h0C000004; // JAL 4 (跳转到地址 4，并将返回地址存入 $31)

        // 测试 J (无条件跳转到 4)
        mem[29] = 32'h08000001; // J 4 (跳转到地址 4)

        // 设置跳转测试寄存器值，确保 J 跳转成功
        mem[30] = 32'h34080001; // ORI $8, $0, 0x01

        // 无条件跳转到 0 号指令
        mem[31] = 32'h08000000; // J 0 (跳转到地址 0)
    end



    assign data = (ce == 1'b1) ? mem[addr[11:2]] : 32'b0; // 地址对齐，非使能输出 0

endmodule
